configuration rtl of try is
    
    
    
end configuration rtl;